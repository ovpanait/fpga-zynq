`timescale 1ns/1ns
`define PERIOD 5

module sha_w_tb();

   // Module instantiation
   reg clk;
   reg reset;
   reg en;
   reg [511:0] M;
   wire [1023:0] W;
   wire en_out;

   sha_w DUT (
		.clk(clk),
		.reset(reset),
		.en(en),
		.M(M),
		.W(W),
		.en_next(en_out)
		);

   // Test setup
   integer     errors;

   // Auxiliary counters
   integer i;

   initial begin
      clk <= 0;
      forever #(`PERIOD) clk = ~clk;
   end

   initial begin
      reset <= 0;
      @(posedge clk); //may need several cycles for reset
      @(negedge clk) reset = 1;
   end

   initial begin
      errors = 0; // reset error count

      // reset inputs to chip
      //chipin1 = 0;
      //chipin2 = 16’ha5;

      // reset simulation parameters
      //resetsim();

      // reset for chip
      //reset_fpga();

      //
      // Add testcases here
      //
`include "test1.sv"

      $display("\nSimulation completed with %d errors\n", errors);
      $stop;
   end

class tester #(int unsigned WIDTH = 32);

   static task verify_output(input [WIDTH-1:0] simulated_value, input [WIDTH-1:0] expected_value);
      begin
	 if (simulated_value[WIDTH-1:0] != expected_value[WIDTH-1:0])
	   begin
	      errors = errors + 1;
	      $display("Simulated Value = %h \n \
	        Expected Value = %h \n \
		errors = %d \n \
		at time = %d\n",
		simulated_value,
		expected_value,
		errors,
		$time);
	   end
end
endtask

endclass

endmodule
