`include "sha.vh"

module sha_block(
	     input 		      clk,
	     input 		      reset,
	     input 		      en,
	     input [`MSG_S-1:0]       M,

	     output [`H_SIZE-1:0] H,
	     output en_next
	     );

wire [`WARR_S-1:0] W[1:0];
wire [`WORD_S-1:0] tmp[7:0];
wire [`WORD_S-1:0] Hin[7:0];
wire en_o[3:0];

localparam K = {
	32'hC67178F2, 32'hBEF9A3F7, 32'hA4506CEB, 32'h90BEFFFA,
	32'h8CC70208, 32'h84C87814, 32'h78A5636F, 32'h748F82EE,
	32'h682E6FF3, 32'h5B9CCA4F, 32'h4ED8AA4A, 32'h391C0CB3,
	32'h34B0BCB5, 32'h2748774C, 32'h1E376C08, 32'h19A4C116,
	32'h106AA070, 32'hF40E3585, 32'hD6990624, 32'hD192E819,
	32'hC76C51A3, 32'hC24B8B70, 32'hA81A664B, 32'hA2BFE8A1,
	32'h92722C85, 32'h81C2C92E, 32'h766A0ABB, 32'h650A7354,
	32'h53380D13, 32'h4D2C6DFC, 32'h2E1B2138, 32'h27B70A85,
	32'h14292967, 32'h06CA6351, 32'hD5A79147, 32'hC6E00BF3,
	32'hBF597FC7, 32'hB00327C8, 32'hA831C66D, 32'h983E5152,
	32'h76F988DA, 32'h5CB0A9DC, 32'h4A7484AA, 32'h2DE92C6F,
	32'h240CA1CC, 32'h0FC19DC6, 32'hEFBE4786, 32'hE49B69C1,
	32'hC19BF174, 32'h9BDC06A7, 32'h80DEB1FE, 32'h72BE5D74,
	32'h550C7DC3, 32'h243185BE, 32'h12835B01, 32'hD807AA98,
	32'hAB1C5ED5, 32'h923F82A4, 32'h59F111F1, 32'h3956C25B,
	32'hE9B5DBA5, 32'hB5C0FBCF, 32'h71374491, 32'h428A2F98
	};


localparam H0 = {
	32'h6a09e667, 32'hbb67ae85, 32'h3c6ef372, 32'ha54ff53a,
	32'h510e527f, 32'h9b05688c, 32'h1f83d9ab, 32'h5be0cd19
	};


// Modules
W_start w_b(
	.clk(clk),
	.reset(reset),
	.en(en),
	.M(M),
	.W(W[0]),
	.en_next(en_o[0]));

W_middle w_e(
	.clk(clk),
	.reset(reset),
	.en(en_o[0]),
	.Win(W[0]),
	.W(W[1]),
	.en_next(en_o[1]));

sha_round round1(
	.clk(clk),
	.reset(reset),
	.en(en_o[1]),

	.a(H0[`VEC_I(7)]),
	.b(H0[`VEC_I(6)]),
	.c(H0[`VEC_I(5)]),
	.d(H0[`VEC_I(4)]),
	.e(H0[`VEC_I(3)]),
	.f(H0[`VEC_I(2)]),
	.g(H0[`VEC_I(1)]),
	.h(H0[`VEC_I(0)]),

	.a_next(tmp[0]),
	.b_next(tmp[1]),
	.c_next(tmp[2]),
	.d_next(tmp[3]),
	.e_next(tmp[4]),
	.f_next(tmp[5]),
	.g_next(tmp[6]),
	.h_next(tmp[7]),

	.K(K[1023:0]),
	.W(W[0]),

	.en_next(en_o[2])
	);

sha_round round2(
	.clk(clk),
	.reset(reset),
	.en(en_o[2]),

	.a(tmp[0]),
	.b(tmp[1]),
	.c(tmp[2]),
	.d(tmp[3]),
	.e(tmp[4]),
	.f(tmp[5]),
	.g(tmp[6]),
	.h(tmp[7]),

	.K(K[2047:1024]),
	.W(W[1]),

	.a_next(Hin[0]),
	.b_next(Hin[1]),
	.c_next(Hin[2]),
	.d_next(Hin[3]),
	.e_next(Hin[4]),
	.f_next(Hin[5]),
	.g_next(Hin[6]),
	.h_next(Hin[7]),

	.en_next(en_o[3])
	);

sha_hash hash_out(
	.clk(clk),
	.reset(reset),
	.en_H(en),
	.en_regs(en_o[3]),

	.H_prev({H0[`VEC_I(7)], H0[`VEC_I(6)], H0[`VEC_I(5)], H0[`VEC_I(4)], H0[`VEC_I(3)], H0[`VEC_I(2)], H0[`VEC_I(1)], H0[`VEC_I(0)]}),
	.a(Hin[0]),
	.b(Hin[1]),
	.c(Hin[2]),
	.d(Hin[3]),
	.e(Hin[4]),
	.f(Hin[5]),
	.g(Hin[6]),
	.h(Hin[7]),

	.H(H),
	.en_o(en_next));

endmodule
